typedef uvm_sequencer#(fifo_tx) wr_sqr;
