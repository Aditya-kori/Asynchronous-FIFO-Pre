typedef uvm_sequencer#(fifo_tx) rd_sqr;
